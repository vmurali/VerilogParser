import Vector::*;
import HaskellLib::*;
import Connectable::*;
import Base::*;
import Primitive::*;
export Types::*;

import RegFile::*;
export RegFile::*;

typedef Bit#(32) VAddr;
typedef Bit#(32) Inst;
typedef Bit#(32) Data;
typedef 32 NumRegs;
typedef TLog#(NumRegs) RegIndexSz;
typedef Bit#(RegIndexSz) RegIndex;
typedef Int#(32) SData;

typedef struct {
  RegIndex index;
  Maybe#(Data) data;
} Wb deriving (Bits, Eq);

typedef union tagged {
  VAddr Load;
  MemWrite Store;
} Mem deriving (Bits, Eq);

typedef struct {
  VAddr pc;
  Bool epoch;
} PcQ deriving (Bits, Eq);

typedef RegFileWrite#(NumRegs, Data) RegWrite;
typedef RegFileWrite#(TExp#(32), Data) MemWrite;

